

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity duck is
    Port (
        v_sync : IN STD_LOGIC;
        pixel_row : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
        pixel_col : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
        bat_x : IN STD_LOGIC_VECTOR (10 DOWNTO 0); -- current bat x position
        bat_y : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
        shoot : IN STD_LOGIC;
        x_position : OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
        y_position : OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
        draw_on : OUT STD_LOGIC;
        X_DIR : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
        hit : OUT STD_LOGIC;
        respawn: IN STD_LOGIC;
        reset: IN STD_LOGIC
     );
end duck;

architecture Behavioral of duck is
    TYPE BUTTON IS (PRESSED,NOT_PRESSED);
    CONSTANT bsize : INTEGER := 8; -- ball size in pixels
    CONSTANT bat_w : INTEGER := 20; -- bat width in pixels
    CONSTANT bat_h : INTEGER := 20; -- bat height in pixels
    -- distance ball moves each frame
    SIGNAL  ball_speed : STD_LOGIC_VECTOR (10 DOWNTO 0) := CONV_STD_LOGIC_VECTOR (2, 11);
    SIGNAL ball_on : STD_LOGIC; -- indicates whether ball is at current pixel position
    SIGNAL game_on : STD_LOGIC := '1'; -- indicates whether ball is in play
    SIGNAL serve : STD_LOGIC := '1';
    SIGNAL nx_hit: STD_LOGIC := '0';
    -- current ball position - intitialized to center of screen
    --SIGNAL ball_x : STD_LOGIC_VECTOR(10 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(400, 11);
    SIGNAL ball_x : STD_LOGIC_VECTOR(10 DOWNTO 0);
    SIGNAL ball_y : STD_LOGIC_VECTOR(10 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(300, 11);
    -- bat vertical position
    --CONSTANT bat_y : STD_LOGIC_VECTOR(10 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(500, 11);
    -- current ball motion - initialized to (+ ball_speed) pixels/frame in both X and Y directions
    SIGNAL ball_x_motion, ball_y_motion : STD_LOGIC_VECTOR(10 DOWNTO 0) := CONV_STD_LOGIC_VECTOR (2, 11);
    SIGNAL shot_state: BUTTON;
    SIGNAL nx_shot_state : BUTTON;
    SIGNAL nx_speed : STD_LOGIC_VECTOR (10 DOWNTO 0);
begin
    x_position <= ball_x;
    y_position <= ball_y;
    draw_on <= game_on;
    
    ck_process : process(v_sync)
    
    begin
    hit <= nx_hit;
    shot_state <= nx_shot_state;
    ball_speed <= nx_speed;
    end process;
    
    
    hitDected : process
    
    BEGIN
    IF reset = '0' THEN
        game_on <= '1';
        nx_speed <= CONV_STD_LOGIC_VECTOR (2, 11);
        ELSE
        IF respawn = '1' THEN
        game_on <= '1';
        nx_hit <= '0';
        ELSE
        WAIT UNTIL rising_edge(v_sync);
        nx_speed <= ball_speed;
        nx_shot_state <= shot_state;
        IF shot_state = NOT_PRESSED THEN
            IF shoot = '1' THEN
                IF (ball_x + bsize/2) >= (bat_x - bat_w) AND
                (ball_x - bsize/2) <= (bat_x + bat_w) AND
                (ball_y + bsize/2) >= (bat_y - bat_h) AND
                (ball_y - bsize/2) <= (bat_y + bat_h) THEN
                    game_on <= '0';
                    nx_hit <= '1';
                    nx_speed <= ball_speed + 1;
                    END IF;
                nx_shot_state <= PRESSED;
            END IF;
        else
            IF shoot = '0' THEN
                nx_shot_state <= NOT_PRESSED;
            ELSE
                nx_shot_state <= PRESSED;
                END IF;
        END IF;
        END IF;
        END IF;
    END PROCESS;
    
    
    mball : PROCESS
        VARIABLE temp : STD_LOGIC_VECTOR (11 DOWNTO 0);
    BEGIN
        WAIT UNTIL rising_edge(v_sync);
        --IF serve = '1' THEN -- test for new serve
          --  ball_x <= X_DIR;
          --  serve <= '0';
           -- game_on <= '1';
           -- ball_y_motion <= (NOT ball_speed) + 1; -- set vspeed to (- ball_speed) pixels

        
        IF ball_y <= bsize THEN -- bounce off top wall
            ball_y_motion <= ball_speed; -- set vspeed to (+ ball_speed) pixels
        ELSIF ball_y + bsize >= 600 THEN -- if ball meets bottom wall
            ball_y_motion <= (NOT ball_speed) + 1; -- set vspeed to (- ball_speed) pixels
            --game_on <= '1'; -- and make ball disappear
        END IF;
        -- allow for bounce off left or right of screen
        IF ball_x + bsize >= 800 THEN -- bounce off right wall
            ball_x_motion <= (NOT ball_speed) + 1; -- set hspeed to (- ball_speed) pixels
        ELSIF ball_x <= bsize THEN -- bounce off left wall
            ball_x_motion <= ball_speed; -- set hspeed to (+ ball_speed) pixels
        END IF;
        -- allow for bounce off bat

        -- compute next ball vertical position
        -- variable temp adds one more bit to calculation to fix unsigned underflow problems
        -- when ball_y is close to zero and ball_y_motion is negative
        temp := ('0' & ball_y) + (ball_y_motion(10) & ball_y_motion);
        IF game_on = '0' THEN
            ball_y <= CONV_STD_LOGIC_VECTOR(799, 11);
            ball_y_motion <= (NOT ball_speed) + 1;
        ELSIF temp(11) = '1' THEN
            ball_y <= (OTHERS => '0');
        ELSE ball_y <= temp(10 DOWNTO 0); -- 9 downto 0
        END IF;
        -- compute next ball horizontal position
        -- variable temp adds one more bit to calculation to fix unsigned underflow problems
        -- when ball_x is close to zero and ball_x_motion is negative
        temp := ('0' & ball_x) + (ball_x_motion(10) & ball_x_motion);
       IF serve = '1' THEN
            ball_x <= x_DIR;
            serve <= '0';
        ELSIF temp(11) = '1' THEN
            ball_x <= (OTHERS => '0');
        ELSE ball_x <= temp(10 DOWNTO 0);
        END IF;
   END PROCESS;
    
end Behavioral;
